lpm_shiftreg16_inst : lpm_shiftreg16 PORT MAP (
		clock	 => clock_sig,
		enable	 => enable_sig,
		shiftin	 => shiftin_sig,
		q	 => q_sig
	);
